/*
 * name: MUX
 * author: btapple
 * description: some multiplexers.
 */

`ifndef __MUX_V__
`define __MUX_V__
`include "./macro.vh"
`timescale 1ns / 1ps

module Mux4 #(parameter WIDTH = 8)
(
    input [WIDTH-1:0] a0,
    input [WIDTH-1:0] a1,
    input [WIDTH-1:0] a2,
    input [WIDTH-1:0] a3,
    input [1:0] select,
    output [WIDTH-1:0] out
);
    assign out= (~(|(select ^ 2'h0)))? a0 :
                (~(|(select ^ 2'h1)))? a1 :
                (~(|(select ^ 2'h2)))? a2 :
                a3;
endmodule // mux4

module Mux2 #(parameter WIDTH = 16)
(
    input [WIDTH-1:0] a0,
    input [WIDTH-1:0] a1,
    input select,
    output [WIDTH-1:0] out
);
    assign out= (~select)?a0:a1;
endmodule // mux2

module Mux3 #(parameter WIDTH = 32)
(
    input [WIDTH-1:0] a0,
    input [WIDTH-1:0] a1,
    input [WIDTH-1:0] a2,
    input [1:0] select,
    output [WIDTH-1:0] out
);
    assign out = (~(|(select ^ 2'h0)))? a0:
                 (~(|(select ^ 2'h1)))? a1:
                 a2;
endmodule // mux3

// module ALUBE_forward_imm_selector(
//     input [`Word] a0,
//     input [`Word] a1,
//     input [`Word] a2,
//     input [`Word] a3,
//     input [1:0] Forward,
//     input Imm,
//     output [`Word] out
// );
//     assign out = (Imm)?a0:
//                  (~(|(Forward ^ `FW_NONEE))) ? a1:
//                  (~(|(Forward ^ `FW_ME)))    ? a2:
//                                                a3;
// endmodule
`endif